** Profile: "SCHEMATIC1-AnalizaBiasPoint"  [ C:\Users\vboxuser\Documents\GitHub\UniRepo\CEA\Lab6MOSFET\Lab6MOSFET-PSpiceFiles\SCHEMATIC1\AnalizaBiasPoint.sim ] 

** Creating circuit file "AnalizaBiasPoint.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OP
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
