** Profile: "SCHEMATIC1-DCSweep_eval"  [ C:\GitHub\UniRepo\CEA\Circuite\test_ex2-PSpiceFiles\SCHEMATIC1\DCSweep_eval.sim ] 

** Creating circuit file "DCSweep_eval.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\mihai\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V2 0 6 0.01 
+ LIN V_V1 0.65 0.73 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
